// $Id: $
// File name:   tb_flex_counter.sv
// Created:     2/2/2018
// Author:      Rochak Chandra
// Lab Section: 337-06
// Version:     1.0  Initial Design Entry
// Description: Test Bench for Flex Counter
